module one_Bit_ADC(
input in1,
input in2,
input vdd,
output out
);
endmodule
