MACRO one_Bit_ADC
  ORIGIN 0 0 ;
  FOREIGN one_Bit_ADC 0 0 ;
  SIZE 11.18 BY 15.12 ;
  PIN OUT
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 7.14 7 8.34 7.28 ;
      LAYER M2 ;
        RECT 8.86 7.84 10.06 8.12 ;
      LAYER M2 ;
        RECT 8.01 7 8.33 7.28 ;
      LAYER M1 ;
        RECT 8.045 7.14 8.295 7.98 ;
      LAYER M2 ;
        RECT 8.17 7.84 9.03 8.12 ;
    END
  END OUT
  PIN VDD
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M3 ;
        RECT 10.18 0.68 10.46 6.88 ;
      LAYER M3 ;
        RECT 10.18 8.24 10.46 14.44 ;
      LAYER M3 ;
        RECT 7.17 8.24 7.45 14.02 ;
      LAYER M3 ;
        RECT 10.18 6.72 10.46 8.4 ;
      LAYER M3 ;
        RECT 10.18 8.635 10.46 9.005 ;
      LAYER M2 ;
        RECT 7.31 8.68 10.32 8.96 ;
      LAYER M3 ;
        RECT 7.17 8.635 7.45 9.005 ;
    END
  END VDD
  PIN IN1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 0.26 10.36 1.46 10.64 ;
    END
  END IN1
  PIN IN2
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 3.7 10.36 4.9 10.64 ;
    END
  END IN2
  OBS 
  LAYER M3 ;
        RECT 4.59 2.78 4.87 7.3 ;
  LAYER M2 ;
        RECT 7.14 2.8 8.34 3.08 ;
  LAYER M3 ;
        RECT 4.59 3.175 4.87 3.545 ;
  LAYER M2 ;
        RECT 4.73 3.22 6.45 3.5 ;
  LAYER M1 ;
        RECT 6.325 2.94 6.575 3.36 ;
  LAYER M2 ;
        RECT 6.45 2.8 7.31 3.08 ;
  LAYER M3 ;
        RECT 9.75 2.78 10.03 7.3 ;
  LAYER M2 ;
        RECT 8.01 2.8 8.33 3.08 ;
  LAYER M3 ;
        RECT 8.03 2.94 8.31 3.36 ;
  LAYER M2 ;
        RECT 8.17 3.22 9.89 3.5 ;
  LAYER M3 ;
        RECT 9.75 3.175 10.03 3.545 ;
  LAYER M2 ;
        RECT 8.01 2.8 8.33 3.08 ;
  LAYER M3 ;
        RECT 8.03 2.78 8.31 3.1 ;
  LAYER M2 ;
        RECT 8.01 3.22 8.33 3.5 ;
  LAYER M3 ;
        RECT 8.03 3.2 8.31 3.52 ;
  LAYER M2 ;
        RECT 9.73 3.22 10.05 3.5 ;
  LAYER M3 ;
        RECT 9.75 3.2 10.03 3.52 ;
  LAYER M2 ;
        RECT 8.01 2.8 8.33 3.08 ;
  LAYER M3 ;
        RECT 8.03 2.78 8.31 3.1 ;
  LAYER M2 ;
        RECT 8.01 3.22 8.33 3.5 ;
  LAYER M3 ;
        RECT 8.03 3.2 8.31 3.52 ;
  LAYER M2 ;
        RECT 9.73 3.22 10.05 3.5 ;
  LAYER M3 ;
        RECT 9.75 3.2 10.03 3.52 ;
  LAYER M2 ;
        RECT 3.7 6.58 4.9 6.86 ;
  LAYER M3 ;
        RECT 3.3 8.24 3.58 14.44 ;
  LAYER M3 ;
        RECT 1.58 8.24 1.86 14.44 ;
  LAYER M2 ;
        RECT 3.44 6.58 3.87 6.86 ;
  LAYER M3 ;
        RECT 3.3 6.72 3.58 8.4 ;
  LAYER M3 ;
        RECT 3.3 9.475 3.58 9.845 ;
  LAYER M2 ;
        RECT 1.72 9.52 3.44 9.8 ;
  LAYER M3 ;
        RECT 1.58 9.475 1.86 9.845 ;
  LAYER M2 ;
        RECT 3.28 6.58 3.6 6.86 ;
  LAYER M3 ;
        RECT 3.3 6.56 3.58 6.88 ;
  LAYER M2 ;
        RECT 3.28 6.58 3.6 6.86 ;
  LAYER M3 ;
        RECT 3.3 6.56 3.58 6.88 ;
  LAYER M2 ;
        RECT 1.56 9.52 1.88 9.8 ;
  LAYER M3 ;
        RECT 1.58 9.5 1.86 9.82 ;
  LAYER M2 ;
        RECT 3.28 6.58 3.6 6.86 ;
  LAYER M3 ;
        RECT 3.3 6.56 3.58 6.88 ;
  LAYER M2 ;
        RECT 3.28 9.52 3.6 9.8 ;
  LAYER M3 ;
        RECT 3.3 9.5 3.58 9.82 ;
  LAYER M2 ;
        RECT 1.56 9.52 1.88 9.8 ;
  LAYER M3 ;
        RECT 1.58 9.5 1.86 9.82 ;
  LAYER M2 ;
        RECT 3.28 6.58 3.6 6.86 ;
  LAYER M3 ;
        RECT 3.3 6.56 3.58 6.88 ;
  LAYER M2 ;
        RECT 3.28 9.52 3.6 9.8 ;
  LAYER M3 ;
        RECT 3.3 9.5 3.58 9.82 ;
  LAYER M3 ;
        RECT 3.73 0.68 4.01 6.46 ;
  LAYER M3 ;
        RECT 6.74 0.68 7.02 6.88 ;
  LAYER M3 ;
        RECT 3.73 3.595 4.01 3.965 ;
  LAYER M2 ;
        RECT 3.87 3.64 6.88 3.92 ;
  LAYER M3 ;
        RECT 6.74 3.595 7.02 3.965 ;
  LAYER M2 ;
        RECT 0.26 14.56 1.46 14.84 ;
  LAYER M3 ;
        RECT 6.31 10.34 6.59 14.86 ;
  LAYER M2 ;
        RECT 1.29 14.56 3.01 14.84 ;
  LAYER M3 ;
        RECT 2.87 13.86 3.15 14.7 ;
  LAYER M4 ;
        RECT 3.01 13.46 6.45 14.26 ;
  LAYER M3 ;
        RECT 6.31 13.675 6.59 14.045 ;
  LAYER M2 ;
        RECT 2.85 14.56 3.17 14.84 ;
  LAYER M3 ;
        RECT 2.87 14.54 3.15 14.86 ;
  LAYER M3 ;
        RECT 2.87 13.675 3.15 14.045 ;
  LAYER M4 ;
        RECT 2.845 13.46 3.175 14.26 ;
  LAYER M3 ;
        RECT 6.31 13.675 6.59 14.045 ;
  LAYER M4 ;
        RECT 6.285 13.46 6.615 14.26 ;
  LAYER M2 ;
        RECT 2.85 14.56 3.17 14.84 ;
  LAYER M3 ;
        RECT 2.87 14.54 3.15 14.86 ;
  LAYER M3 ;
        RECT 2.87 13.675 3.15 14.045 ;
  LAYER M4 ;
        RECT 2.845 13.46 3.175 14.26 ;
  LAYER M3 ;
        RECT 6.31 13.675 6.59 14.045 ;
  LAYER M4 ;
        RECT 6.285 13.46 6.615 14.26 ;
  LAYER M2 ;
        RECT 3.7 14.56 4.9 14.84 ;
  LAYER M2 ;
        RECT 6.28 14.14 7.48 14.42 ;
  LAYER M2 ;
        RECT 8.86 12.04 10.06 12.32 ;
  LAYER M2 ;
        RECT 4.57 14.56 4.89 14.84 ;
  LAYER M1 ;
        RECT 4.605 14.7 4.855 15.12 ;
  LAYER M2 ;
        RECT 4.73 14.98 6.02 15.26 ;
  LAYER M3 ;
        RECT 5.88 14.28 6.16 15.12 ;
  LAYER M2 ;
        RECT 6.02 14.14 6.45 14.42 ;
  LAYER M2 ;
        RECT 7.31 14.14 7.74 14.42 ;
  LAYER M3 ;
        RECT 7.6 12.18 7.88 14.28 ;
  LAYER M2 ;
        RECT 7.74 12.04 9.03 12.32 ;
  LAYER M1 ;
        RECT 4.605 14.615 4.855 14.785 ;
  LAYER M2 ;
        RECT 4.56 14.56 4.9 14.84 ;
  LAYER M1 ;
        RECT 4.605 15.035 4.855 15.205 ;
  LAYER M2 ;
        RECT 4.56 14.98 4.9 15.26 ;
  LAYER M2 ;
        RECT 5.86 14.14 6.18 14.42 ;
  LAYER M3 ;
        RECT 5.88 14.12 6.16 14.44 ;
  LAYER M2 ;
        RECT 5.86 14.98 6.18 15.26 ;
  LAYER M3 ;
        RECT 5.88 14.96 6.16 15.28 ;
  LAYER M1 ;
        RECT 4.605 14.615 4.855 14.785 ;
  LAYER M2 ;
        RECT 4.56 14.56 4.9 14.84 ;
  LAYER M1 ;
        RECT 4.605 15.035 4.855 15.205 ;
  LAYER M2 ;
        RECT 4.56 14.98 4.9 15.26 ;
  LAYER M2 ;
        RECT 5.86 14.14 6.18 14.42 ;
  LAYER M3 ;
        RECT 5.88 14.12 6.16 14.44 ;
  LAYER M2 ;
        RECT 5.86 14.98 6.18 15.26 ;
  LAYER M3 ;
        RECT 5.88 14.96 6.16 15.28 ;
  LAYER M1 ;
        RECT 4.605 14.615 4.855 14.785 ;
  LAYER M2 ;
        RECT 4.56 14.56 4.9 14.84 ;
  LAYER M1 ;
        RECT 4.605 15.035 4.855 15.205 ;
  LAYER M2 ;
        RECT 4.56 14.98 4.9 15.26 ;
  LAYER M2 ;
        RECT 5.86 14.14 6.18 14.42 ;
  LAYER M3 ;
        RECT 5.88 14.12 6.16 14.44 ;
  LAYER M2 ;
        RECT 5.86 14.98 6.18 15.26 ;
  LAYER M3 ;
        RECT 5.88 14.96 6.16 15.28 ;
  LAYER M2 ;
        RECT 7.58 12.04 7.9 12.32 ;
  LAYER M3 ;
        RECT 7.6 12.02 7.88 12.34 ;
  LAYER M2 ;
        RECT 7.58 14.14 7.9 14.42 ;
  LAYER M3 ;
        RECT 7.6 14.12 7.88 14.44 ;
  LAYER M1 ;
        RECT 4.605 14.615 4.855 14.785 ;
  LAYER M2 ;
        RECT 4.56 14.56 4.9 14.84 ;
  LAYER M1 ;
        RECT 4.605 15.035 4.855 15.205 ;
  LAYER M2 ;
        RECT 4.56 14.98 4.9 15.26 ;
  LAYER M2 ;
        RECT 5.86 14.14 6.18 14.42 ;
  LAYER M3 ;
        RECT 5.88 14.12 6.16 14.44 ;
  LAYER M2 ;
        RECT 5.86 14.98 6.18 15.26 ;
  LAYER M3 ;
        RECT 5.88 14.96 6.16 15.28 ;
  LAYER M2 ;
        RECT 7.58 12.04 7.9 12.32 ;
  LAYER M3 ;
        RECT 7.6 12.02 7.88 12.34 ;
  LAYER M2 ;
        RECT 7.58 14.14 7.9 14.42 ;
  LAYER M3 ;
        RECT 7.6 14.12 7.88 14.44 ;
  LAYER M1 ;
        RECT 4.605 3.695 4.855 7.225 ;
  LAYER M1 ;
        RECT 4.605 2.435 4.855 3.445 ;
  LAYER M1 ;
        RECT 4.605 0.335 4.855 1.345 ;
  LAYER M1 ;
        RECT 5.035 3.695 5.285 7.225 ;
  LAYER M1 ;
        RECT 4.175 3.695 4.425 7.225 ;
  LAYER M1 ;
        RECT 3.745 3.695 3.995 7.225 ;
  LAYER M1 ;
        RECT 3.745 2.435 3.995 3.445 ;
  LAYER M1 ;
        RECT 3.745 0.335 3.995 1.345 ;
  LAYER M1 ;
        RECT 3.315 3.695 3.565 7.225 ;
  LAYER M2 ;
        RECT 3.7 2.8 4.9 3.08 ;
  LAYER M2 ;
        RECT 4.56 7 5.76 7.28 ;
  LAYER M2 ;
        RECT 3.27 6.16 5.33 6.44 ;
  LAYER M2 ;
        RECT 3.7 0.7 4.9 0.98 ;
  LAYER M3 ;
        RECT 4.59 2.78 4.87 7.3 ;
  LAYER M2 ;
        RECT 3.7 6.58 4.9 6.86 ;
  LAYER M3 ;
        RECT 3.73 0.68 4.01 6.46 ;
  LAYER M1 ;
        RECT 7.185 3.695 7.435 7.225 ;
  LAYER M1 ;
        RECT 7.185 2.435 7.435 3.445 ;
  LAYER M1 ;
        RECT 7.185 0.335 7.435 1.345 ;
  LAYER M1 ;
        RECT 7.615 3.695 7.865 7.225 ;
  LAYER M1 ;
        RECT 6.755 3.695 7.005 7.225 ;
  LAYER M2 ;
        RECT 6.71 6.58 7.91 6.86 ;
  LAYER M2 ;
        RECT 6.71 0.7 7.91 0.98 ;
  LAYER M2 ;
        RECT 7.14 7 8.34 7.28 ;
  LAYER M2 ;
        RECT 7.14 2.8 8.34 3.08 ;
  LAYER M3 ;
        RECT 6.74 0.68 7.02 6.88 ;
  LAYER M1 ;
        RECT 6.325 11.255 6.575 14.785 ;
  LAYER M1 ;
        RECT 6.325 9.995 6.575 11.005 ;
  LAYER M1 ;
        RECT 6.325 7.895 6.575 8.905 ;
  LAYER M1 ;
        RECT 5.895 11.255 6.145 14.785 ;
  LAYER M1 ;
        RECT 6.755 11.255 7.005 14.785 ;
  LAYER M1 ;
        RECT 7.185 11.255 7.435 14.785 ;
  LAYER M1 ;
        RECT 7.185 9.995 7.435 11.005 ;
  LAYER M1 ;
        RECT 7.185 7.895 7.435 8.905 ;
  LAYER M1 ;
        RECT 7.615 11.255 7.865 14.785 ;
  LAYER M2 ;
        RECT 6.28 10.36 7.48 10.64 ;
  LAYER M2 ;
        RECT 5.42 14.56 6.62 14.84 ;
  LAYER M2 ;
        RECT 5.85 13.72 7.91 14 ;
  LAYER M2 ;
        RECT 6.28 8.26 7.48 8.54 ;
  LAYER M3 ;
        RECT 6.31 10.34 6.59 14.86 ;
  LAYER M2 ;
        RECT 6.28 14.14 7.48 14.42 ;
  LAYER M3 ;
        RECT 7.17 8.24 7.45 14.02 ;
  LAYER M1 ;
        RECT 9.765 3.695 10.015 7.225 ;
  LAYER M1 ;
        RECT 9.765 2.435 10.015 3.445 ;
  LAYER M1 ;
        RECT 9.765 0.335 10.015 1.345 ;
  LAYER M1 ;
        RECT 9.335 3.695 9.585 7.225 ;
  LAYER M1 ;
        RECT 10.195 3.695 10.445 7.225 ;
  LAYER M2 ;
        RECT 8.86 2.8 10.06 3.08 ;
  LAYER M2 ;
        RECT 8.86 7 10.06 7.28 ;
  LAYER M2 ;
        RECT 9.29 6.58 10.49 6.86 ;
  LAYER M2 ;
        RECT 9.29 0.7 10.49 0.98 ;
  LAYER M3 ;
        RECT 9.75 2.78 10.03 7.3 ;
  LAYER M3 ;
        RECT 10.18 0.68 10.46 6.88 ;
  LAYER M1 ;
        RECT 1.165 11.255 1.415 14.785 ;
  LAYER M1 ;
        RECT 1.165 9.995 1.415 11.005 ;
  LAYER M1 ;
        RECT 1.165 7.895 1.415 8.905 ;
  LAYER M1 ;
        RECT 0.735 11.255 0.985 14.785 ;
  LAYER M1 ;
        RECT 1.595 11.255 1.845 14.785 ;
  LAYER M2 ;
        RECT 0.69 14.14 1.89 14.42 ;
  LAYER M2 ;
        RECT 0.69 8.26 1.89 8.54 ;
  LAYER M2 ;
        RECT 0.26 14.56 1.46 14.84 ;
  LAYER M2 ;
        RECT 0.26 10.36 1.46 10.64 ;
  LAYER M3 ;
        RECT 1.58 8.24 1.86 14.44 ;
  LAYER M1 ;
        RECT 3.745 11.255 3.995 14.785 ;
  LAYER M1 ;
        RECT 3.745 9.995 3.995 11.005 ;
  LAYER M1 ;
        RECT 3.745 7.895 3.995 8.905 ;
  LAYER M1 ;
        RECT 4.175 11.255 4.425 14.785 ;
  LAYER M1 ;
        RECT 3.315 11.255 3.565 14.785 ;
  LAYER M2 ;
        RECT 3.27 14.14 4.47 14.42 ;
  LAYER M2 ;
        RECT 3.27 8.26 4.47 8.54 ;
  LAYER M2 ;
        RECT 3.7 14.56 4.9 14.84 ;
  LAYER M2 ;
        RECT 3.7 10.36 4.9 10.64 ;
  LAYER M3 ;
        RECT 3.3 8.24 3.58 14.44 ;
  LAYER M1 ;
        RECT 9.765 7.895 10.015 11.425 ;
  LAYER M1 ;
        RECT 9.765 11.675 10.015 12.685 ;
  LAYER M1 ;
        RECT 9.765 13.775 10.015 14.785 ;
  LAYER M1 ;
        RECT 9.335 7.895 9.585 11.425 ;
  LAYER M1 ;
        RECT 10.195 7.895 10.445 11.425 ;
  LAYER M2 ;
        RECT 9.29 8.26 10.49 8.54 ;
  LAYER M2 ;
        RECT 9.29 14.14 10.49 14.42 ;
  LAYER M2 ;
        RECT 8.86 7.84 10.06 8.12 ;
  LAYER M2 ;
        RECT 8.86 12.04 10.06 12.32 ;
  LAYER M3 ;
        RECT 10.18 8.24 10.46 14.44 ;
  END 
END one_Bit_ADC
