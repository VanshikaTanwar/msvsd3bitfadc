VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO Ring_Osc_Analog
  CLASS BLOCK ;
  FOREIGN Ring_Osc_Analog ;
  ORIGIN 0.000 -0.150 ;
  SIZE 5.160 BY 29.940 ;
  OBS
      LAYER pwell ;
        RECT 2.365 28.710 2.795 30.090 ;
        RECT 1.895 24.860 3.265 26.170 ;
      LAYER nwell ;
        RECT 1.290 15.120 3.870 22.680 ;
        RECT 0.000 7.560 5.160 15.120 ;
      LAYER pwell ;
        RECT 0.605 4.070 1.975 5.380 ;
        RECT 3.185 4.070 4.555 5.380 ;
        RECT 1.075 0.150 1.505 1.530 ;
        RECT 3.655 0.150 4.085 1.530 ;
      LAYER li1 ;
        RECT 2.455 28.895 2.705 29.905 ;
        RECT 2.455 26.795 2.705 27.805 ;
        RECT 2.025 23.015 2.275 26.545 ;
        RECT 2.455 23.015 2.705 26.545 ;
        RECT 2.885 23.015 3.135 26.545 ;
        RECT 2.025 18.815 2.275 22.345 ;
        RECT 2.455 18.815 2.705 22.345 ;
        RECT 2.885 18.815 3.135 22.345 ;
        RECT 1.165 13.775 1.415 14.785 ;
        RECT 1.165 11.675 1.415 12.685 ;
        RECT 0.735 7.895 0.985 11.425 ;
        RECT 1.165 7.895 1.415 11.425 ;
        RECT 1.595 7.895 1.845 11.425 ;
        RECT 2.025 7.895 2.275 18.145 ;
        RECT 2.455 17.555 2.705 18.565 ;
        RECT 3.315 17.975 3.565 27.385 ;
        RECT 2.455 15.455 2.705 16.465 ;
        RECT 3.745 13.775 3.995 14.785 ;
        RECT 0.735 3.695 0.985 7.225 ;
        RECT 1.165 3.695 1.415 7.225 ;
        RECT 1.595 3.695 1.845 7.225 ;
        RECT 1.165 2.435 1.415 3.445 ;
        RECT 2.455 2.855 2.705 12.265 ;
        RECT 3.745 11.675 3.995 12.685 ;
        RECT 3.315 7.895 3.565 11.425 ;
        RECT 3.745 7.895 3.995 11.425 ;
        RECT 4.175 7.895 4.425 11.425 ;
        RECT 3.315 3.695 3.565 7.225 ;
        RECT 3.745 3.695 3.995 7.225 ;
        RECT 4.175 3.695 4.425 7.225 ;
        RECT 3.745 2.435 3.995 3.445 ;
        RECT 1.165 0.335 1.415 1.345 ;
        RECT 3.745 0.335 3.995 1.345 ;
      LAYER mcon ;
        RECT 2.495 29.315 2.665 29.485 ;
        RECT 2.495 27.215 2.665 27.385 ;
        RECT 3.355 27.215 3.525 27.385 ;
        RECT 2.065 23.435 2.235 23.605 ;
        RECT 2.495 23.015 2.665 23.185 ;
        RECT 2.925 23.435 3.095 23.605 ;
        RECT 2.065 21.755 2.235 21.925 ;
        RECT 2.495 22.175 2.665 22.345 ;
        RECT 2.925 21.755 3.095 21.925 ;
        RECT 2.065 17.975 2.235 18.145 ;
        RECT 1.205 14.195 1.375 14.365 ;
        RECT 1.205 12.095 1.375 12.265 ;
        RECT 0.775 8.315 0.945 8.485 ;
        RECT 1.205 7.895 1.375 8.065 ;
        RECT 1.635 8.315 1.805 8.485 ;
        RECT 2.495 17.975 2.665 18.145 ;
        RECT 3.355 17.975 3.525 18.145 ;
        RECT 2.495 15.875 2.665 16.045 ;
        RECT 3.785 14.195 3.955 14.365 ;
        RECT 2.065 7.895 2.235 8.065 ;
        RECT 2.495 12.095 2.665 12.265 ;
        RECT 3.785 12.095 3.955 12.265 ;
        RECT 3.355 8.315 3.525 8.485 ;
        RECT 3.785 7.895 3.955 8.065 ;
        RECT 4.215 8.315 4.385 8.485 ;
        RECT 0.775 6.635 0.945 6.805 ;
        RECT 1.205 7.055 1.375 7.225 ;
        RECT 1.635 6.635 1.805 6.805 ;
        RECT 2.495 7.055 2.665 7.225 ;
        RECT 1.205 2.855 1.375 3.025 ;
        RECT 3.355 6.635 3.525 6.805 ;
        RECT 3.785 7.055 3.955 7.225 ;
        RECT 4.215 6.635 4.385 6.805 ;
        RECT 2.495 2.855 2.665 3.025 ;
        RECT 3.785 2.855 3.955 3.025 ;
        RECT 1.205 0.755 1.375 0.925 ;
        RECT 3.785 0.755 3.955 0.925 ;
      LAYER met1 ;
        RECT 1.980 29.260 3.180 29.540 ;
        RECT 2.410 27.160 3.610 27.440 ;
        RECT 1.980 23.380 3.180 23.660 ;
        RECT 2.410 22.960 3.610 23.240 ;
        RECT 2.410 22.120 4.030 22.400 ;
        RECT 1.980 21.700 3.180 21.980 ;
        RECT 1.980 17.920 3.610 18.200 ;
        RECT 1.980 15.820 3.180 16.100 ;
        RECT 1.990 14.560 3.600 14.840 ;
        RECT 0.690 14.140 1.890 14.420 ;
        RECT 3.270 14.140 4.470 14.420 ;
        RECT 0.260 12.040 2.750 12.320 ;
        RECT 3.700 12.040 4.900 12.320 ;
        RECT 1.560 11.200 3.600 11.480 ;
        RECT 0.690 8.260 1.890 8.540 ;
        RECT 3.270 8.260 4.470 8.540 ;
        RECT 0.260 7.840 2.320 8.120 ;
        RECT 3.700 7.840 4.900 8.120 ;
        RECT 0.260 7.000 1.460 7.280 ;
        RECT 2.410 7.000 4.900 7.280 ;
        RECT 0.690 6.580 1.890 6.860 ;
        RECT 3.270 6.580 4.470 6.860 ;
        RECT 1.560 3.640 3.600 3.920 ;
        RECT 0.260 2.800 2.750 3.080 ;
        RECT 3.700 2.800 4.900 3.080 ;
        RECT 0.690 0.700 1.890 0.980 ;
        RECT 3.270 0.700 4.470 0.980 ;
      LAYER via ;
        RECT 2.020 29.270 2.280 29.530 ;
        RECT 2.020 23.390 2.280 23.650 ;
        RECT 2.880 22.970 3.140 23.230 ;
        RECT 2.880 22.130 3.140 22.390 ;
        RECT 3.740 22.130 4.000 22.390 ;
        RECT 2.020 21.710 2.280 21.970 ;
        RECT 2.020 15.830 2.280 16.090 ;
        RECT 2.020 14.570 2.280 14.830 ;
        RECT 3.310 14.570 3.570 14.830 ;
        RECT 1.590 14.150 1.850 14.410 ;
        RECT 3.310 14.150 3.570 14.410 ;
        RECT 3.740 12.050 4.000 12.310 ;
        RECT 4.170 12.050 4.430 12.310 ;
        RECT 1.590 11.210 1.850 11.470 ;
        RECT 3.310 11.210 3.570 11.470 ;
        RECT 1.590 8.270 1.850 8.530 ;
        RECT 3.310 8.270 3.570 8.530 ;
        RECT 0.730 7.850 0.990 8.110 ;
        RECT 3.740 7.850 4.000 8.110 ;
        RECT 0.730 7.010 0.990 7.270 ;
        RECT 3.740 7.010 4.000 7.270 ;
        RECT 1.590 6.590 1.850 6.850 ;
        RECT 3.310 6.590 3.570 6.850 ;
        RECT 1.590 3.650 1.850 3.910 ;
        RECT 3.310 3.650 3.570 3.910 ;
        RECT 4.170 2.810 4.430 3.070 ;
        RECT 1.590 0.710 1.850 0.970 ;
        RECT 3.310 0.710 3.570 0.970 ;
      LAYER met2 ;
        RECT 2.010 22.495 2.290 29.560 ;
        RECT 2.870 22.100 3.150 23.260 ;
        RECT 2.010 14.540 2.290 22.000 ;
        RECT 1.580 8.240 1.860 14.440 ;
        RECT 3.300 8.240 3.580 14.860 ;
        RECT 3.730 12.020 4.010 22.420 ;
        RECT 0.720 6.980 1.000 8.140 ;
        RECT 1.580 0.680 1.860 7.745 ;
        RECT 3.730 6.980 4.010 8.140 ;
        RECT 3.300 0.680 3.580 6.880 ;
        RECT 4.160 2.780 4.440 12.340 ;
      LAYER via2 ;
        RECT 2.010 22.540 2.290 22.820 ;
        RECT 1.580 7.420 1.860 7.700 ;
      LAYER met3 ;
        RECT 1.315 22.280 2.315 23.080 ;
        RECT 1.315 7.160 1.885 7.960 ;
      LAYER via3 ;
        RECT 1.320 22.520 1.640 22.840 ;
        RECT 1.320 7.400 1.640 7.720 ;
      LAYER met4 ;
        RECT 0.890 7.395 2.070 22.845 ;
  END
END Ring_Osc_Analog
END LIBRARY

