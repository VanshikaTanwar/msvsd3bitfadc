module Ring_Osc_Analog (
 output Vout
 );
endmodule
